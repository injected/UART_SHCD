----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    10:48:20 11/13/2010 
-- Design Name: 
-- Module Name:    ARMADEUS_DUMMY - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity E_ARMADEUS_DUMMY is
	Port 
	( 
		E_ARMADEUS_DUMMY_Reset: 				IN  STD_LOGIC;
		E_ARMADEUS_DUMMY_Clock_In:					IN  STD_LOGIC
);
end E_ARMADEUS_DUMMY;

architecture ARMADEUS_DUMMY_A of E_ARMADEUS_DUMMY is

begin


end ARMADEUS_DUMMY_A;

